-- SQ_GEN.VHD (a peripheral module for SCOMP)
-- 2020.10.10
--
-- Generates a square wave with period dependant on value
-- sent from SCOMP.

LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.numeric_std.ALL;
USE LPM.LPM_COMPONENTS.ALL;


ENTITY SQ_GEN IS
	PORT(
		CLOCK, -- 100 kHz clock
		RESETN,
		CS       : IN STD_LOGIC;
		IO_DATA  : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		IO_WRITE : IN    STD_LOGIC;
		SQ       : OUT STD_LOGIC;
		DURATION_EN : IN STD_LOGIC;
		SPACE_EN: IN STD_LOGIC;
		PAUSE_EN: IN STD_LOGIC
	);
END SQ_GEN;


ARCHITECTURE a OF SQ_GEN IS
	constant clock_freq : INTEGER := 100000;
	constant half_freq : INTEGER := clock_freq/2; -- 50% duty cycle
	
	SIGNAL COUNT : INTEGER RANGE 0 to 10000;
	SIGNAL D        : STD_LOGIC;
	SIGNAL ENABLED : STD_LOGIC;
	
	SIGNAL PAUSED : STD_LOGIC;
	
	SIGNAL COMPARE : INTEGER RANGE 0 to 10000;
	signal next_compare : integer range 0 to 10000;
	
	signal duration_cycles : integer;
	signal next_duration_cycles : integer;
	
	signal inputs_started : integer;
	signal inputs_accepted : integer;
	signal has_space : std_logic;
	
	SIGNAL TICKER : INTEGER RANGE 0 to clock_freq/8; -- 8 Hz rollover. 16 Hz is too fast.
	signal duration_cycle_counter : integer;
	
	type to_comp_map is array (0 to 2093) of integer;
	constant mapping : to_comp_map := (
		0,
		half_freq/1,
		half_freq/2,
		half_freq/3,
		half_freq/4,
		half_freq/5,
		half_freq/6,
		half_freq/7,
		half_freq/8,
		half_freq/9,
		half_freq/10,
		half_freq/11,
		half_freq/12,
		half_freq/13,
		half_freq/14,
		half_freq/15,
		half_freq/16,
		half_freq/17,
		half_freq/18,
		half_freq/19,
		half_freq/20,
		half_freq/21,
		half_freq/22,
		half_freq/23,
		half_freq/24,
		half_freq/25,
		half_freq/26,
		half_freq/27,
		half_freq/28,
		half_freq/29,
		half_freq/30,
		half_freq/31,
		half_freq/32,
		half_freq/33,
		half_freq/34,
		half_freq/35,
		half_freq/36,
		half_freq/37,
		half_freq/38,
		half_freq/39,
		half_freq/40,
		half_freq/41,
		half_freq/42,
		half_freq/43,
		half_freq/44,
		half_freq/45,
		half_freq/46,
		half_freq/47,
		half_freq/48,
		half_freq/49,
		half_freq/50,
		half_freq/51,
		half_freq/52,
		half_freq/53,
		half_freq/54,
		half_freq/55,
		half_freq/56,
		half_freq/57,
		half_freq/58,
		half_freq/59,
		half_freq/60,
		half_freq/61,
		half_freq/62,
		half_freq/63,
		half_freq/64,
		half_freq/65,
		half_freq/66,
		half_freq/67,
		half_freq/68,
		half_freq/69,
		half_freq/70,
		half_freq/71,
		half_freq/72,
		half_freq/73,
		half_freq/74,
		half_freq/75,
		half_freq/76,
		half_freq/77,
		half_freq/78,
		half_freq/79,
		half_freq/80,
		half_freq/81,
		half_freq/82,
		half_freq/83,
		half_freq/84,
		half_freq/85,
		half_freq/86,
		half_freq/87,
		half_freq/88,
		half_freq/89,
		half_freq/90,
		half_freq/91,
		half_freq/92,
		half_freq/93,
		half_freq/94,
		half_freq/95,
		half_freq/96,
		half_freq/97,
		half_freq/98,
		half_freq/99,
		half_freq/100,
		half_freq/101,
		half_freq/102,
		half_freq/103,
		half_freq/104,
		half_freq/105,
		half_freq/106,
		half_freq/107,
		half_freq/108,
		half_freq/109,
		half_freq/110,
		half_freq/111,
		half_freq/112,
		half_freq/113,
		half_freq/114,
		half_freq/115,
		half_freq/116,
		half_freq/117,
		half_freq/118,
		half_freq/119,
		half_freq/120,
		half_freq/121,
		half_freq/122,
		half_freq/123,
		half_freq/124,
		half_freq/125,
		half_freq/126,
		half_freq/127,
		half_freq/128,
		half_freq/129,
		half_freq/130,
		half_freq/131,
		half_freq/132,
		half_freq/133,
		half_freq/134,
		half_freq/135,
		half_freq/136,
		half_freq/137,
		half_freq/138,
		half_freq/139,
		half_freq/140,
		half_freq/141,
		half_freq/142,
		half_freq/143,
		half_freq/144,
		half_freq/145,
		half_freq/146,
		half_freq/147,
		half_freq/148,
		half_freq/149,
		half_freq/150,
		half_freq/151,
		half_freq/152,
		half_freq/153,
		half_freq/154,
		half_freq/155,
		half_freq/156,
		half_freq/157,
		half_freq/158,
		half_freq/159,
		half_freq/160,
		half_freq/161,
		half_freq/162,
		half_freq/163,
		half_freq/164,
		half_freq/165,
		half_freq/166,
		half_freq/167,
		half_freq/168,
		half_freq/169,
		half_freq/170,
		half_freq/171,
		half_freq/172,
		half_freq/173,
		half_freq/174,
		half_freq/175,
		half_freq/176,
		half_freq/177,
		half_freq/178,
		half_freq/179,
		half_freq/180,
		half_freq/181,
		half_freq/182,
		half_freq/183,
		half_freq/184,
		half_freq/185,
		half_freq/186,
		half_freq/187,
		half_freq/188,
		half_freq/189,
		half_freq/190,
		half_freq/191,
		half_freq/192,
		half_freq/193,
		half_freq/194,
		half_freq/195,
		half_freq/196,
		half_freq/197,
		half_freq/198,
		half_freq/199,
		half_freq/200,
		half_freq/201,
		half_freq/202,
		half_freq/203,
		half_freq/204,
		half_freq/205,
		half_freq/206,
		half_freq/207,
		half_freq/208,
		half_freq/209,
		half_freq/210,
		half_freq/211,
		half_freq/212,
		half_freq/213,
		half_freq/214,
		half_freq/215,
		half_freq/216,
		half_freq/217,
		half_freq/218,
		half_freq/219,
		half_freq/220,
		half_freq/221,
		half_freq/222,
		half_freq/223,
		half_freq/224,
		half_freq/225,
		half_freq/226,
		half_freq/227,
		half_freq/228,
		half_freq/229,
		half_freq/230,
		half_freq/231,
		half_freq/232,
		half_freq/233,
		half_freq/234,
		half_freq/235,
		half_freq/236,
		half_freq/237,
		half_freq/238,
		half_freq/239,
		half_freq/240,
		half_freq/241,
		half_freq/242,
		half_freq/243,
		half_freq/244,
		half_freq/245,
		half_freq/246,
		half_freq/247,
		half_freq/248,
		half_freq/249,
		half_freq/250,
		half_freq/251,
		half_freq/252,
		half_freq/253,
		half_freq/254,
		half_freq/255,
		half_freq/256,
		half_freq/257,
		half_freq/258,
		half_freq/259,
		half_freq/260,
		half_freq/261,
		half_freq/262,
		half_freq/263,
		half_freq/264,
		half_freq/265,
		half_freq/266,
		half_freq/267,
		half_freq/268,
		half_freq/269,
		half_freq/270,
		half_freq/271,
		half_freq/272,
		half_freq/273,
		half_freq/274,
		half_freq/275,
		half_freq/276,
		half_freq/277,
		half_freq/278,
		half_freq/279,
		half_freq/280,
		half_freq/281,
		half_freq/282,
		half_freq/283,
		half_freq/284,
		half_freq/285,
		half_freq/286,
		half_freq/287,
		half_freq/288,
		half_freq/289,
		half_freq/290,
		half_freq/291,
		half_freq/292,
		half_freq/293,
		half_freq/294,
		half_freq/295,
		half_freq/296,
		half_freq/297,
		half_freq/298,
		half_freq/299,
		half_freq/300,
		half_freq/301,
		half_freq/302,
		half_freq/303,
		half_freq/304,
		half_freq/305,
		half_freq/306,
		half_freq/307,
		half_freq/308,
		half_freq/309,
		half_freq/310,
		half_freq/311,
		half_freq/312,
		half_freq/313,
		half_freq/314,
		half_freq/315,
		half_freq/316,
		half_freq/317,
		half_freq/318,
		half_freq/319,
		half_freq/320,
		half_freq/321,
		half_freq/322,
		half_freq/323,
		half_freq/324,
		half_freq/325,
		half_freq/326,
		half_freq/327,
		half_freq/328,
		half_freq/329,
		half_freq/330,
		half_freq/331,
		half_freq/332,
		half_freq/333,
		half_freq/334,
		half_freq/335,
		half_freq/336,
		half_freq/337,
		half_freq/338,
		half_freq/339,
		half_freq/340,
		half_freq/341,
		half_freq/342,
		half_freq/343,
		half_freq/344,
		half_freq/345,
		half_freq/346,
		half_freq/347,
		half_freq/348,
		half_freq/349,
		half_freq/350,
		half_freq/351,
		half_freq/352,
		half_freq/353,
		half_freq/354,
		half_freq/355,
		half_freq/356,
		half_freq/357,
		half_freq/358,
		half_freq/359,
		half_freq/360,
		half_freq/361,
		half_freq/362,
		half_freq/363,
		half_freq/364,
		half_freq/365,
		half_freq/366,
		half_freq/367,
		half_freq/368,
		half_freq/369,
		half_freq/370,
		half_freq/371,
		half_freq/372,
		half_freq/373,
		half_freq/374,
		half_freq/375,
		half_freq/376,
		half_freq/377,
		half_freq/378,
		half_freq/379,
		half_freq/380,
		half_freq/381,
		half_freq/382,
		half_freq/383,
		half_freq/384,
		half_freq/385,
		half_freq/386,
		half_freq/387,
		half_freq/388,
		half_freq/389,
		half_freq/390,
		half_freq/391,
		half_freq/392,
		half_freq/393,
		half_freq/394,
		half_freq/395,
		half_freq/396,
		half_freq/397,
		half_freq/398,
		half_freq/399,
		half_freq/400,
		half_freq/401,
		half_freq/402,
		half_freq/403,
		half_freq/404,
		half_freq/405,
		half_freq/406,
		half_freq/407,
		half_freq/408,
		half_freq/409,
		half_freq/410,
		half_freq/411,
		half_freq/412,
		half_freq/413,
		half_freq/414,
		half_freq/415,
		half_freq/416,
		half_freq/417,
		half_freq/418,
		half_freq/419,
		half_freq/420,
		half_freq/421,
		half_freq/422,
		half_freq/423,
		half_freq/424,
		half_freq/425,
		half_freq/426,
		half_freq/427,
		half_freq/428,
		half_freq/429,
		half_freq/430,
		half_freq/431,
		half_freq/432,
		half_freq/433,
		half_freq/434,
		half_freq/435,
		half_freq/436,
		half_freq/437,
		half_freq/438,
		half_freq/439,
		half_freq/440,
		half_freq/441,
		half_freq/442,
		half_freq/443,
		half_freq/444,
		half_freq/445,
		half_freq/446,
		half_freq/447,
		half_freq/448,
		half_freq/449,
		half_freq/450,
		half_freq/451,
		half_freq/452,
		half_freq/453,
		half_freq/454,
		half_freq/455,
		half_freq/456,
		half_freq/457,
		half_freq/458,
		half_freq/459,
		half_freq/460,
		half_freq/461,
		half_freq/462,
		half_freq/463,
		half_freq/464,
		half_freq/465,
		half_freq/466,
		half_freq/467,
		half_freq/468,
		half_freq/469,
		half_freq/470,
		half_freq/471,
		half_freq/472,
		half_freq/473,
		half_freq/474,
		half_freq/475,
		half_freq/476,
		half_freq/477,
		half_freq/478,
		half_freq/479,
		half_freq/480,
		half_freq/481,
		half_freq/482,
		half_freq/483,
		half_freq/484,
		half_freq/485,
		half_freq/486,
		half_freq/487,
		half_freq/488,
		half_freq/489,
		half_freq/490,
		half_freq/491,
		half_freq/492,
		half_freq/493,
		half_freq/494,
		half_freq/495,
		half_freq/496,
		half_freq/497,
		half_freq/498,
		half_freq/499,
		half_freq/500,
		half_freq/501,
		half_freq/502,
		half_freq/503,
		half_freq/504,
		half_freq/505,
		half_freq/506,
		half_freq/507,
		half_freq/508,
		half_freq/509,
		half_freq/510,
		half_freq/511,
		half_freq/512,
		half_freq/513,
		half_freq/514,
		half_freq/515,
		half_freq/516,
		half_freq/517,
		half_freq/518,
		half_freq/519,
		half_freq/520,
		half_freq/521,
		half_freq/522,
		half_freq/523,
		half_freq/524,
		half_freq/525,
		half_freq/526,
		half_freq/527,
		half_freq/528,
		half_freq/529,
		half_freq/530,
		half_freq/531,
		half_freq/532,
		half_freq/533,
		half_freq/534,
		half_freq/535,
		half_freq/536,
		half_freq/537,
		half_freq/538,
		half_freq/539,
		half_freq/540,
		half_freq/541,
		half_freq/542,
		half_freq/543,
		half_freq/544,
		half_freq/545,
		half_freq/546,
		half_freq/547,
		half_freq/548,
		half_freq/549,
		half_freq/550,
		half_freq/551,
		half_freq/552,
		half_freq/553,
		half_freq/554,
		half_freq/555,
		half_freq/556,
		half_freq/557,
		half_freq/558,
		half_freq/559,
		half_freq/560,
		half_freq/561,
		half_freq/562,
		half_freq/563,
		half_freq/564,
		half_freq/565,
		half_freq/566,
		half_freq/567,
		half_freq/568,
		half_freq/569,
		half_freq/570,
		half_freq/571,
		half_freq/572,
		half_freq/573,
		half_freq/574,
		half_freq/575,
		half_freq/576,
		half_freq/577,
		half_freq/578,
		half_freq/579,
		half_freq/580,
		half_freq/581,
		half_freq/582,
		half_freq/583,
		half_freq/584,
		half_freq/585,
		half_freq/586,
		half_freq/587,
		half_freq/588,
		half_freq/589,
		half_freq/590,
		half_freq/591,
		half_freq/592,
		half_freq/593,
		half_freq/594,
		half_freq/595,
		half_freq/596,
		half_freq/597,
		half_freq/598,
		half_freq/599,
		half_freq/600,
		half_freq/601,
		half_freq/602,
		half_freq/603,
		half_freq/604,
		half_freq/605,
		half_freq/606,
		half_freq/607,
		half_freq/608,
		half_freq/609,
		half_freq/610,
		half_freq/611,
		half_freq/612,
		half_freq/613,
		half_freq/614,
		half_freq/615,
		half_freq/616,
		half_freq/617,
		half_freq/618,
		half_freq/619,
		half_freq/620,
		half_freq/621,
		half_freq/622,
		half_freq/623,
		half_freq/624,
		half_freq/625,
		half_freq/626,
		half_freq/627,
		half_freq/628,
		half_freq/629,
		half_freq/630,
		half_freq/631,
		half_freq/632,
		half_freq/633,
		half_freq/634,
		half_freq/635,
		half_freq/636,
		half_freq/637,
		half_freq/638,
		half_freq/639,
		half_freq/640,
		half_freq/641,
		half_freq/642,
		half_freq/643,
		half_freq/644,
		half_freq/645,
		half_freq/646,
		half_freq/647,
		half_freq/648,
		half_freq/649,
		half_freq/650,
		half_freq/651,
		half_freq/652,
		half_freq/653,
		half_freq/654,
		half_freq/655,
		half_freq/656,
		half_freq/657,
		half_freq/658,
		half_freq/659,
		half_freq/660,
		half_freq/661,
		half_freq/662,
		half_freq/663,
		half_freq/664,
		half_freq/665,
		half_freq/666,
		half_freq/667,
		half_freq/668,
		half_freq/669,
		half_freq/670,
		half_freq/671,
		half_freq/672,
		half_freq/673,
		half_freq/674,
		half_freq/675,
		half_freq/676,
		half_freq/677,
		half_freq/678,
		half_freq/679,
		half_freq/680,
		half_freq/681,
		half_freq/682,
		half_freq/683,
		half_freq/684,
		half_freq/685,
		half_freq/686,
		half_freq/687,
		half_freq/688,
		half_freq/689,
		half_freq/690,
		half_freq/691,
		half_freq/692,
		half_freq/693,
		half_freq/694,
		half_freq/695,
		half_freq/696,
		half_freq/697,
		half_freq/698,
		half_freq/699,
		half_freq/700,
		half_freq/701,
		half_freq/702,
		half_freq/703,
		half_freq/704,
		half_freq/705,
		half_freq/706,
		half_freq/707,
		half_freq/708,
		half_freq/709,
		half_freq/710,
		half_freq/711,
		half_freq/712,
		half_freq/713,
		half_freq/714,
		half_freq/715,
		half_freq/716,
		half_freq/717,
		half_freq/718,
		half_freq/719,
		half_freq/720,
		half_freq/721,
		half_freq/722,
		half_freq/723,
		half_freq/724,
		half_freq/725,
		half_freq/726,
		half_freq/727,
		half_freq/728,
		half_freq/729,
		half_freq/730,
		half_freq/731,
		half_freq/732,
		half_freq/733,
		half_freq/734,
		half_freq/735,
		half_freq/736,
		half_freq/737,
		half_freq/738,
		half_freq/739,
		half_freq/740,
		half_freq/741,
		half_freq/742,
		half_freq/743,
		half_freq/744,
		half_freq/745,
		half_freq/746,
		half_freq/747,
		half_freq/748,
		half_freq/749,
		half_freq/750,
		half_freq/751,
		half_freq/752,
		half_freq/753,
		half_freq/754,
		half_freq/755,
		half_freq/756,
		half_freq/757,
		half_freq/758,
		half_freq/759,
		half_freq/760,
		half_freq/761,
		half_freq/762,
		half_freq/763,
		half_freq/764,
		half_freq/765,
		half_freq/766,
		half_freq/767,
		half_freq/768,
		half_freq/769,
		half_freq/770,
		half_freq/771,
		half_freq/772,
		half_freq/773,
		half_freq/774,
		half_freq/775,
		half_freq/776,
		half_freq/777,
		half_freq/778,
		half_freq/779,
		half_freq/780,
		half_freq/781,
		half_freq/782,
		half_freq/783,
		half_freq/784,
		half_freq/785,
		half_freq/786,
		half_freq/787,
		half_freq/788,
		half_freq/789,
		half_freq/790,
		half_freq/791,
		half_freq/792,
		half_freq/793,
		half_freq/794,
		half_freq/795,
		half_freq/796,
		half_freq/797,
		half_freq/798,
		half_freq/799,
		half_freq/800,
		half_freq/801,
		half_freq/802,
		half_freq/803,
		half_freq/804,
		half_freq/805,
		half_freq/806,
		half_freq/807,
		half_freq/808,
		half_freq/809,
		half_freq/810,
		half_freq/811,
		half_freq/812,
		half_freq/813,
		half_freq/814,
		half_freq/815,
		half_freq/816,
		half_freq/817,
		half_freq/818,
		half_freq/819,
		half_freq/820,
		half_freq/821,
		half_freq/822,
		half_freq/823,
		half_freq/824,
		half_freq/825,
		half_freq/826,
		half_freq/827,
		half_freq/828,
		half_freq/829,
		half_freq/830,
		half_freq/831,
		half_freq/832,
		half_freq/833,
		half_freq/834,
		half_freq/835,
		half_freq/836,
		half_freq/837,
		half_freq/838,
		half_freq/839,
		half_freq/840,
		half_freq/841,
		half_freq/842,
		half_freq/843,
		half_freq/844,
		half_freq/845,
		half_freq/846,
		half_freq/847,
		half_freq/848,
		half_freq/849,
		half_freq/850,
		half_freq/851,
		half_freq/852,
		half_freq/853,
		half_freq/854,
		half_freq/855,
		half_freq/856,
		half_freq/857,
		half_freq/858,
		half_freq/859,
		half_freq/860,
		half_freq/861,
		half_freq/862,
		half_freq/863,
		half_freq/864,
		half_freq/865,
		half_freq/866,
		half_freq/867,
		half_freq/868,
		half_freq/869,
		half_freq/870,
		half_freq/871,
		half_freq/872,
		half_freq/873,
		half_freq/874,
		half_freq/875,
		half_freq/876,
		half_freq/877,
		half_freq/878,
		half_freq/879,
		half_freq/880,
		half_freq/881,
		half_freq/882,
		half_freq/883,
		half_freq/884,
		half_freq/885,
		half_freq/886,
		half_freq/887,
		half_freq/888,
		half_freq/889,
		half_freq/890,
		half_freq/891,
		half_freq/892,
		half_freq/893,
		half_freq/894,
		half_freq/895,
		half_freq/896,
		half_freq/897,
		half_freq/898,
		half_freq/899,
		half_freq/900,
		half_freq/901,
		half_freq/902,
		half_freq/903,
		half_freq/904,
		half_freq/905,
		half_freq/906,
		half_freq/907,
		half_freq/908,
		half_freq/909,
		half_freq/910,
		half_freq/911,
		half_freq/912,
		half_freq/913,
		half_freq/914,
		half_freq/915,
		half_freq/916,
		half_freq/917,
		half_freq/918,
		half_freq/919,
		half_freq/920,
		half_freq/921,
		half_freq/922,
		half_freq/923,
		half_freq/924,
		half_freq/925,
		half_freq/926,
		half_freq/927,
		half_freq/928,
		half_freq/929,
		half_freq/930,
		half_freq/931,
		half_freq/932,
		half_freq/933,
		half_freq/934,
		half_freq/935,
		half_freq/936,
		half_freq/937,
		half_freq/938,
		half_freq/939,
		half_freq/940,
		half_freq/941,
		half_freq/942,
		half_freq/943,
		half_freq/944,
		half_freq/945,
		half_freq/946,
		half_freq/947,
		half_freq/948,
		half_freq/949,
		half_freq/950,
		half_freq/951,
		half_freq/952,
		half_freq/953,
		half_freq/954,
		half_freq/955,
		half_freq/956,
		half_freq/957,
		half_freq/958,
		half_freq/959,
		half_freq/960,
		half_freq/961,
		half_freq/962,
		half_freq/963,
		half_freq/964,
		half_freq/965,
		half_freq/966,
		half_freq/967,
		half_freq/968,
		half_freq/969,
		half_freq/970,
		half_freq/971,
		half_freq/972,
		half_freq/973,
		half_freq/974,
		half_freq/975,
		half_freq/976,
		half_freq/977,
		half_freq/978,
		half_freq/979,
		half_freq/980,
		half_freq/981,
		half_freq/982,
		half_freq/983,
		half_freq/984,
		half_freq/985,
		half_freq/986,
		half_freq/987,
		half_freq/988,
		half_freq/989,
		half_freq/990,
		half_freq/991,
		half_freq/992,
		half_freq/993,
		half_freq/994,
		half_freq/995,
		half_freq/996,
		half_freq/997,
		half_freq/998,
		half_freq/999,
		half_freq/1000,
		half_freq/1001,
		half_freq/1002,
		half_freq/1003,
		half_freq/1004,
		half_freq/1005,
		half_freq/1006,
		half_freq/1007,
		half_freq/1008,
		half_freq/1009,
		half_freq/1010,
		half_freq/1011,
		half_freq/1012,
		half_freq/1013,
		half_freq/1014,
		half_freq/1015,
		half_freq/1016,
		half_freq/1017,
		half_freq/1018,
		half_freq/1019,
		half_freq/1020,
		half_freq/1021,
		half_freq/1022,
		half_freq/1023,
		half_freq/1024,
		half_freq/1025,
		half_freq/1026,
		half_freq/1027,
		half_freq/1028,
		half_freq/1029,
		half_freq/1030,
		half_freq/1031,
		half_freq/1032,
		half_freq/1033,
		half_freq/1034,
		half_freq/1035,
		half_freq/1036,
		half_freq/1037,
		half_freq/1038,
		half_freq/1039,
		half_freq/1040,
		half_freq/1041,
		half_freq/1042,
		half_freq/1043,
		half_freq/1044,
		half_freq/1045,
		half_freq/1046,
		half_freq/1047,
		half_freq/1048,
		half_freq/1049,
		half_freq/1050,
		half_freq/1051,
		half_freq/1052,
		half_freq/1053,
		half_freq/1054,
		half_freq/1055,
		half_freq/1056,
		half_freq/1057,
		half_freq/1058,
		half_freq/1059,
		half_freq/1060,
		half_freq/1061,
		half_freq/1062,
		half_freq/1063,
		half_freq/1064,
		half_freq/1065,
		half_freq/1066,
		half_freq/1067,
		half_freq/1068,
		half_freq/1069,
		half_freq/1070,
		half_freq/1071,
		half_freq/1072,
		half_freq/1073,
		half_freq/1074,
		half_freq/1075,
		half_freq/1076,
		half_freq/1077,
		half_freq/1078,
		half_freq/1079,
		half_freq/1080,
		half_freq/1081,
		half_freq/1082,
		half_freq/1083,
		half_freq/1084,
		half_freq/1085,
		half_freq/1086,
		half_freq/1087,
		half_freq/1088,
		half_freq/1089,
		half_freq/1090,
		half_freq/1091,
		half_freq/1092,
		half_freq/1093,
		half_freq/1094,
		half_freq/1095,
		half_freq/1096,
		half_freq/1097,
		half_freq/1098,
		half_freq/1099,
		half_freq/1100,
		half_freq/1101,
		half_freq/1102,
		half_freq/1103,
		half_freq/1104,
		half_freq/1105,
		half_freq/1106,
		half_freq/1107,
		half_freq/1108,
		half_freq/1109,
		half_freq/1110,
		half_freq/1111,
		half_freq/1112,
		half_freq/1113,
		half_freq/1114,
		half_freq/1115,
		half_freq/1116,
		half_freq/1117,
		half_freq/1118,
		half_freq/1119,
		half_freq/1120,
		half_freq/1121,
		half_freq/1122,
		half_freq/1123,
		half_freq/1124,
		half_freq/1125,
		half_freq/1126,
		half_freq/1127,
		half_freq/1128,
		half_freq/1129,
		half_freq/1130,
		half_freq/1131,
		half_freq/1132,
		half_freq/1133,
		half_freq/1134,
		half_freq/1135,
		half_freq/1136,
		half_freq/1137,
		half_freq/1138,
		half_freq/1139,
		half_freq/1140,
		half_freq/1141,
		half_freq/1142,
		half_freq/1143,
		half_freq/1144,
		half_freq/1145,
		half_freq/1146,
		half_freq/1147,
		half_freq/1148,
		half_freq/1149,
		half_freq/1150,
		half_freq/1151,
		half_freq/1152,
		half_freq/1153,
		half_freq/1154,
		half_freq/1155,
		half_freq/1156,
		half_freq/1157,
		half_freq/1158,
		half_freq/1159,
		half_freq/1160,
		half_freq/1161,
		half_freq/1162,
		half_freq/1163,
		half_freq/1164,
		half_freq/1165,
		half_freq/1166,
		half_freq/1167,
		half_freq/1168,
		half_freq/1169,
		half_freq/1170,
		half_freq/1171,
		half_freq/1172,
		half_freq/1173,
		half_freq/1174,
		half_freq/1175,
		half_freq/1176,
		half_freq/1177,
		half_freq/1178,
		half_freq/1179,
		half_freq/1180,
		half_freq/1181,
		half_freq/1182,
		half_freq/1183,
		half_freq/1184,
		half_freq/1185,
		half_freq/1186,
		half_freq/1187,
		half_freq/1188,
		half_freq/1189,
		half_freq/1190,
		half_freq/1191,
		half_freq/1192,
		half_freq/1193,
		half_freq/1194,
		half_freq/1195,
		half_freq/1196,
		half_freq/1197,
		half_freq/1198,
		half_freq/1199,
		half_freq/1200,
		half_freq/1201,
		half_freq/1202,
		half_freq/1203,
		half_freq/1204,
		half_freq/1205,
		half_freq/1206,
		half_freq/1207,
		half_freq/1208,
		half_freq/1209,
		half_freq/1210,
		half_freq/1211,
		half_freq/1212,
		half_freq/1213,
		half_freq/1214,
		half_freq/1215,
		half_freq/1216,
		half_freq/1217,
		half_freq/1218,
		half_freq/1219,
		half_freq/1220,
		half_freq/1221,
		half_freq/1222,
		half_freq/1223,
		half_freq/1224,
		half_freq/1225,
		half_freq/1226,
		half_freq/1227,
		half_freq/1228,
		half_freq/1229,
		half_freq/1230,
		half_freq/1231,
		half_freq/1232,
		half_freq/1233,
		half_freq/1234,
		half_freq/1235,
		half_freq/1236,
		half_freq/1237,
		half_freq/1238,
		half_freq/1239,
		half_freq/1240,
		half_freq/1241,
		half_freq/1242,
		half_freq/1243,
		half_freq/1244,
		half_freq/1245,
		half_freq/1246,
		half_freq/1247,
		half_freq/1248,
		half_freq/1249,
		half_freq/1250,
		half_freq/1251,
		half_freq/1252,
		half_freq/1253,
		half_freq/1254,
		half_freq/1255,
		half_freq/1256,
		half_freq/1257,
		half_freq/1258,
		half_freq/1259,
		half_freq/1260,
		half_freq/1261,
		half_freq/1262,
		half_freq/1263,
		half_freq/1264,
		half_freq/1265,
		half_freq/1266,
		half_freq/1267,
		half_freq/1268,
		half_freq/1269,
		half_freq/1270,
		half_freq/1271,
		half_freq/1272,
		half_freq/1273,
		half_freq/1274,
		half_freq/1275,
		half_freq/1276,
		half_freq/1277,
		half_freq/1278,
		half_freq/1279,
		half_freq/1280,
		half_freq/1281,
		half_freq/1282,
		half_freq/1283,
		half_freq/1284,
		half_freq/1285,
		half_freq/1286,
		half_freq/1287,
		half_freq/1288,
		half_freq/1289,
		half_freq/1290,
		half_freq/1291,
		half_freq/1292,
		half_freq/1293,
		half_freq/1294,
		half_freq/1295,
		half_freq/1296,
		half_freq/1297,
		half_freq/1298,
		half_freq/1299,
		half_freq/1300,
		half_freq/1301,
		half_freq/1302,
		half_freq/1303,
		half_freq/1304,
		half_freq/1305,
		half_freq/1306,
		half_freq/1307,
		half_freq/1308,
		half_freq/1309,
		half_freq/1310,
		half_freq/1311,
		half_freq/1312,
		half_freq/1313,
		half_freq/1314,
		half_freq/1315,
		half_freq/1316,
		half_freq/1317,
		half_freq/1318,
		half_freq/1319,
		half_freq/1320,
		half_freq/1321,
		half_freq/1322,
		half_freq/1323,
		half_freq/1324,
		half_freq/1325,
		half_freq/1326,
		half_freq/1327,
		half_freq/1328,
		half_freq/1329,
		half_freq/1330,
		half_freq/1331,
		half_freq/1332,
		half_freq/1333,
		half_freq/1334,
		half_freq/1335,
		half_freq/1336,
		half_freq/1337,
		half_freq/1338,
		half_freq/1339,
		half_freq/1340,
		half_freq/1341,
		half_freq/1342,
		half_freq/1343,
		half_freq/1344,
		half_freq/1345,
		half_freq/1346,
		half_freq/1347,
		half_freq/1348,
		half_freq/1349,
		half_freq/1350,
		half_freq/1351,
		half_freq/1352,
		half_freq/1353,
		half_freq/1354,
		half_freq/1355,
		half_freq/1356,
		half_freq/1357,
		half_freq/1358,
		half_freq/1359,
		half_freq/1360,
		half_freq/1361,
		half_freq/1362,
		half_freq/1363,
		half_freq/1364,
		half_freq/1365,
		half_freq/1366,
		half_freq/1367,
		half_freq/1368,
		half_freq/1369,
		half_freq/1370,
		half_freq/1371,
		half_freq/1372,
		half_freq/1373,
		half_freq/1374,
		half_freq/1375,
		half_freq/1376,
		half_freq/1377,
		half_freq/1378,
		half_freq/1379,
		half_freq/1380,
		half_freq/1381,
		half_freq/1382,
		half_freq/1383,
		half_freq/1384,
		half_freq/1385,
		half_freq/1386,
		half_freq/1387,
		half_freq/1388,
		half_freq/1389,
		half_freq/1390,
		half_freq/1391,
		half_freq/1392,
		half_freq/1393,
		half_freq/1394,
		half_freq/1395,
		half_freq/1396,
		half_freq/1397,
		half_freq/1398,
		half_freq/1399,
		half_freq/1400,
		half_freq/1401,
		half_freq/1402,
		half_freq/1403,
		half_freq/1404,
		half_freq/1405,
		half_freq/1406,
		half_freq/1407,
		half_freq/1408,
		half_freq/1409,
		half_freq/1410,
		half_freq/1411,
		half_freq/1412,
		half_freq/1413,
		half_freq/1414,
		half_freq/1415,
		half_freq/1416,
		half_freq/1417,
		half_freq/1418,
		half_freq/1419,
		half_freq/1420,
		half_freq/1421,
		half_freq/1422,
		half_freq/1423,
		half_freq/1424,
		half_freq/1425,
		half_freq/1426,
		half_freq/1427,
		half_freq/1428,
		half_freq/1429,
		half_freq/1430,
		half_freq/1431,
		half_freq/1432,
		half_freq/1433,
		half_freq/1434,
		half_freq/1435,
		half_freq/1436,
		half_freq/1437,
		half_freq/1438,
		half_freq/1439,
		half_freq/1440,
		half_freq/1441,
		half_freq/1442,
		half_freq/1443,
		half_freq/1444,
		half_freq/1445,
		half_freq/1446,
		half_freq/1447,
		half_freq/1448,
		half_freq/1449,
		half_freq/1450,
		half_freq/1451,
		half_freq/1452,
		half_freq/1453,
		half_freq/1454,
		half_freq/1455,
		half_freq/1456,
		half_freq/1457,
		half_freq/1458,
		half_freq/1459,
		half_freq/1460,
		half_freq/1461,
		half_freq/1462,
		half_freq/1463,
		half_freq/1464,
		half_freq/1465,
		half_freq/1466,
		half_freq/1467,
		half_freq/1468,
		half_freq/1469,
		half_freq/1470,
		half_freq/1471,
		half_freq/1472,
		half_freq/1473,
		half_freq/1474,
		half_freq/1475,
		half_freq/1476,
		half_freq/1477,
		half_freq/1478,
		half_freq/1479,
		half_freq/1480,
		half_freq/1481,
		half_freq/1482,
		half_freq/1483,
		half_freq/1484,
		half_freq/1485,
		half_freq/1486,
		half_freq/1487,
		half_freq/1488,
		half_freq/1489,
		half_freq/1490,
		half_freq/1491,
		half_freq/1492,
		half_freq/1493,
		half_freq/1494,
		half_freq/1495,
		half_freq/1496,
		half_freq/1497,
		half_freq/1498,
		half_freq/1499,
		half_freq/1500,
		half_freq/1501,
		half_freq/1502,
		half_freq/1503,
		half_freq/1504,
		half_freq/1505,
		half_freq/1506,
		half_freq/1507,
		half_freq/1508,
		half_freq/1509,
		half_freq/1510,
		half_freq/1511,
		half_freq/1512,
		half_freq/1513,
		half_freq/1514,
		half_freq/1515,
		half_freq/1516,
		half_freq/1517,
		half_freq/1518,
		half_freq/1519,
		half_freq/1520,
		half_freq/1521,
		half_freq/1522,
		half_freq/1523,
		half_freq/1524,
		half_freq/1525,
		half_freq/1526,
		half_freq/1527,
		half_freq/1528,
		half_freq/1529,
		half_freq/1530,
		half_freq/1531,
		half_freq/1532,
		half_freq/1533,
		half_freq/1534,
		half_freq/1535,
		half_freq/1536,
		half_freq/1537,
		half_freq/1538,
		half_freq/1539,
		half_freq/1540,
		half_freq/1541,
		half_freq/1542,
		half_freq/1543,
		half_freq/1544,
		half_freq/1545,
		half_freq/1546,
		half_freq/1547,
		half_freq/1548,
		half_freq/1549,
		half_freq/1550,
		half_freq/1551,
		half_freq/1552,
		half_freq/1553,
		half_freq/1554,
		half_freq/1555,
		half_freq/1556,
		half_freq/1557,
		half_freq/1558,
		half_freq/1559,
		half_freq/1560,
		half_freq/1561,
		half_freq/1562,
		half_freq/1563,
		half_freq/1564,
		half_freq/1565,
		half_freq/1566,
		half_freq/1567,
		half_freq/1568,
		half_freq/1569,
		half_freq/1570,
		half_freq/1571,
		half_freq/1572,
		half_freq/1573,
		half_freq/1574,
		half_freq/1575,
		half_freq/1576,
		half_freq/1577,
		half_freq/1578,
		half_freq/1579,
		half_freq/1580,
		half_freq/1581,
		half_freq/1582,
		half_freq/1583,
		half_freq/1584,
		half_freq/1585,
		half_freq/1586,
		half_freq/1587,
		half_freq/1588,
		half_freq/1589,
		half_freq/1590,
		half_freq/1591,
		half_freq/1592,
		half_freq/1593,
		half_freq/1594,
		half_freq/1595,
		half_freq/1596,
		half_freq/1597,
		half_freq/1598,
		half_freq/1599,
		half_freq/1600,
		half_freq/1601,
		half_freq/1602,
		half_freq/1603,
		half_freq/1604,
		half_freq/1605,
		half_freq/1606,
		half_freq/1607,
		half_freq/1608,
		half_freq/1609,
		half_freq/1610,
		half_freq/1611,
		half_freq/1612,
		half_freq/1613,
		half_freq/1614,
		half_freq/1615,
		half_freq/1616,
		half_freq/1617,
		half_freq/1618,
		half_freq/1619,
		half_freq/1620,
		half_freq/1621,
		half_freq/1622,
		half_freq/1623,
		half_freq/1624,
		half_freq/1625,
		half_freq/1626,
		half_freq/1627,
		half_freq/1628,
		half_freq/1629,
		half_freq/1630,
		half_freq/1631,
		half_freq/1632,
		half_freq/1633,
		half_freq/1634,
		half_freq/1635,
		half_freq/1636,
		half_freq/1637,
		half_freq/1638,
		half_freq/1639,
		half_freq/1640,
		half_freq/1641,
		half_freq/1642,
		half_freq/1643,
		half_freq/1644,
		half_freq/1645,
		half_freq/1646,
		half_freq/1647,
		half_freq/1648,
		half_freq/1649,
		half_freq/1650,
		half_freq/1651,
		half_freq/1652,
		half_freq/1653,
		half_freq/1654,
		half_freq/1655,
		half_freq/1656,
		half_freq/1657,
		half_freq/1658,
		half_freq/1659,
		half_freq/1660,
		half_freq/1661,
		half_freq/1662,
		half_freq/1663,
		half_freq/1664,
		half_freq/1665,
		half_freq/1666,
		half_freq/1667,
		half_freq/1668,
		half_freq/1669,
		half_freq/1670,
		half_freq/1671,
		half_freq/1672,
		half_freq/1673,
		half_freq/1674,
		half_freq/1675,
		half_freq/1676,
		half_freq/1677,
		half_freq/1678,
		half_freq/1679,
		half_freq/1680,
		half_freq/1681,
		half_freq/1682,
		half_freq/1683,
		half_freq/1684,
		half_freq/1685,
		half_freq/1686,
		half_freq/1687,
		half_freq/1688,
		half_freq/1689,
		half_freq/1690,
		half_freq/1691,
		half_freq/1692,
		half_freq/1693,
		half_freq/1694,
		half_freq/1695,
		half_freq/1696,
		half_freq/1697,
		half_freq/1698,
		half_freq/1699,
		half_freq/1700,
		half_freq/1701,
		half_freq/1702,
		half_freq/1703,
		half_freq/1704,
		half_freq/1705,
		half_freq/1706,
		half_freq/1707,
		half_freq/1708,
		half_freq/1709,
		half_freq/1710,
		half_freq/1711,
		half_freq/1712,
		half_freq/1713,
		half_freq/1714,
		half_freq/1715,
		half_freq/1716,
		half_freq/1717,
		half_freq/1718,
		half_freq/1719,
		half_freq/1720,
		half_freq/1721,
		half_freq/1722,
		half_freq/1723,
		half_freq/1724,
		half_freq/1725,
		half_freq/1726,
		half_freq/1727,
		half_freq/1728,
		half_freq/1729,
		half_freq/1730,
		half_freq/1731,
		half_freq/1732,
		half_freq/1733,
		half_freq/1734,
		half_freq/1735,
		half_freq/1736,
		half_freq/1737,
		half_freq/1738,
		half_freq/1739,
		half_freq/1740,
		half_freq/1741,
		half_freq/1742,
		half_freq/1743,
		half_freq/1744,
		half_freq/1745,
		half_freq/1746,
		half_freq/1747,
		half_freq/1748,
		half_freq/1749,
		half_freq/1750,
		half_freq/1751,
		half_freq/1752,
		half_freq/1753,
		half_freq/1754,
		half_freq/1755,
		half_freq/1756,
		half_freq/1757,
		half_freq/1758,
		half_freq/1759,
		half_freq/1760,
		half_freq/1761,
		half_freq/1762,
		half_freq/1763,
		half_freq/1764,
		half_freq/1765,
		half_freq/1766,
		half_freq/1767,
		half_freq/1768,
		half_freq/1769,
		half_freq/1770,
		half_freq/1771,
		half_freq/1772,
		half_freq/1773,
		half_freq/1774,
		half_freq/1775,
		half_freq/1776,
		half_freq/1777,
		half_freq/1778,
		half_freq/1779,
		half_freq/1780,
		half_freq/1781,
		half_freq/1782,
		half_freq/1783,
		half_freq/1784,
		half_freq/1785,
		half_freq/1786,
		half_freq/1787,
		half_freq/1788,
		half_freq/1789,
		half_freq/1790,
		half_freq/1791,
		half_freq/1792,
		half_freq/1793,
		half_freq/1794,
		half_freq/1795,
		half_freq/1796,
		half_freq/1797,
		half_freq/1798,
		half_freq/1799,
		half_freq/1800,
		half_freq/1801,
		half_freq/1802,
		half_freq/1803,
		half_freq/1804,
		half_freq/1805,
		half_freq/1806,
		half_freq/1807,
		half_freq/1808,
		half_freq/1809,
		half_freq/1810,
		half_freq/1811,
		half_freq/1812,
		half_freq/1813,
		half_freq/1814,
		half_freq/1815,
		half_freq/1816,
		half_freq/1817,
		half_freq/1818,
		half_freq/1819,
		half_freq/1820,
		half_freq/1821,
		half_freq/1822,
		half_freq/1823,
		half_freq/1824,
		half_freq/1825,
		half_freq/1826,
		half_freq/1827,
		half_freq/1828,
		half_freq/1829,
		half_freq/1830,
		half_freq/1831,
		half_freq/1832,
		half_freq/1833,
		half_freq/1834,
		half_freq/1835,
		half_freq/1836,
		half_freq/1837,
		half_freq/1838,
		half_freq/1839,
		half_freq/1840,
		half_freq/1841,
		half_freq/1842,
		half_freq/1843,
		half_freq/1844,
		half_freq/1845,
		half_freq/1846,
		half_freq/1847,
		half_freq/1848,
		half_freq/1849,
		half_freq/1850,
		half_freq/1851,
		half_freq/1852,
		half_freq/1853,
		half_freq/1854,
		half_freq/1855,
		half_freq/1856,
		half_freq/1857,
		half_freq/1858,
		half_freq/1859,
		half_freq/1860,
		half_freq/1861,
		half_freq/1862,
		half_freq/1863,
		half_freq/1864,
		half_freq/1865,
		half_freq/1866,
		half_freq/1867,
		half_freq/1868,
		half_freq/1869,
		half_freq/1870,
		half_freq/1871,
		half_freq/1872,
		half_freq/1873,
		half_freq/1874,
		half_freq/1875,
		half_freq/1876,
		half_freq/1877,
		half_freq/1878,
		half_freq/1879,
		half_freq/1880,
		half_freq/1881,
		half_freq/1882,
		half_freq/1883,
		half_freq/1884,
		half_freq/1885,
		half_freq/1886,
		half_freq/1887,
		half_freq/1888,
		half_freq/1889,
		half_freq/1890,
		half_freq/1891,
		half_freq/1892,
		half_freq/1893,
		half_freq/1894,
		half_freq/1895,
		half_freq/1896,
		half_freq/1897,
		half_freq/1898,
		half_freq/1899,
		half_freq/1900,
		half_freq/1901,
		half_freq/1902,
		half_freq/1903,
		half_freq/1904,
		half_freq/1905,
		half_freq/1906,
		half_freq/1907,
		half_freq/1908,
		half_freq/1909,
		half_freq/1910,
		half_freq/1911,
		half_freq/1912,
		half_freq/1913,
		half_freq/1914,
		half_freq/1915,
		half_freq/1916,
		half_freq/1917,
		half_freq/1918,
		half_freq/1919,
		half_freq/1920,
		half_freq/1921,
		half_freq/1922,
		half_freq/1923,
		half_freq/1924,
		half_freq/1925,
		half_freq/1926,
		half_freq/1927,
		half_freq/1928,
		half_freq/1929,
		half_freq/1930,
		half_freq/1931,
		half_freq/1932,
		half_freq/1933,
		half_freq/1934,
		half_freq/1935,
		half_freq/1936,
		half_freq/1937,
		half_freq/1938,
		half_freq/1939,
		half_freq/1940,
		half_freq/1941,
		half_freq/1942,
		half_freq/1943,
		half_freq/1944,
		half_freq/1945,
		half_freq/1946,
		half_freq/1947,
		half_freq/1948,
		half_freq/1949,
		half_freq/1950,
		half_freq/1951,
		half_freq/1952,
		half_freq/1953,
		half_freq/1954,
		half_freq/1955,
		half_freq/1956,
		half_freq/1957,
		half_freq/1958,
		half_freq/1959,
		half_freq/1960,
		half_freq/1961,
		half_freq/1962,
		half_freq/1963,
		half_freq/1964,
		half_freq/1965,
		half_freq/1966,
		half_freq/1967,
		half_freq/1968,
		half_freq/1969,
		half_freq/1970,
		half_freq/1971,
		half_freq/1972,
		half_freq/1973,
		half_freq/1974,
		half_freq/1975,
		half_freq/1976,
		half_freq/1977,
		half_freq/1978,
		half_freq/1979,
		half_freq/1980,
		half_freq/1981,
		half_freq/1982,
		half_freq/1983,
		half_freq/1984,
		half_freq/1985,
		half_freq/1986,
		half_freq/1987,
		half_freq/1988,
		half_freq/1989,
		half_freq/1990,
		half_freq/1991,
		half_freq/1992,
		half_freq/1993,
		half_freq/1994,
		half_freq/1995,
		half_freq/1996,
		half_freq/1997,
		half_freq/1998,
		half_freq/1999,
		half_freq/2000,
		half_freq/2001,
		half_freq/2002,
		half_freq/2003,
		half_freq/2004,
		half_freq/2005,
		half_freq/2006,
		half_freq/2007,
		half_freq/2008,
		half_freq/2009,
		half_freq/2010,
		half_freq/2011,
		half_freq/2012,
		half_freq/2013,
		half_freq/2014,
		half_freq/2015,
		half_freq/2016,
		half_freq/2017,
		half_freq/2018,
		half_freq/2019,
		half_freq/2020,
		half_freq/2021,
		half_freq/2022,
		half_freq/2023,
		half_freq/2024,
		half_freq/2025,
		half_freq/2026,
		half_freq/2027,
		half_freq/2028,
		half_freq/2029,
		half_freq/2030,
		half_freq/2031,
		half_freq/2032,
		half_freq/2033,
		half_freq/2034,
		half_freq/2035,
		half_freq/2036,
		half_freq/2037,
		half_freq/2038,
		half_freq/2039,
		half_freq/2040,
		half_freq/2041,
		half_freq/2042,
		half_freq/2043,
		half_freq/2044,
		half_freq/2045,
		half_freq/2046,
		half_freq/2047,
		half_freq/2048,
		half_freq/2049,
		half_freq/2050,
		half_freq/2051,
		half_freq/2052,
		half_freq/2053,
		half_freq/2054,
		half_freq/2055,
		half_freq/2056,
		half_freq/2057,
		half_freq/2058,
		half_freq/2059,
		half_freq/2060,
		half_freq/2061,
		half_freq/2062,
		half_freq/2063,
		half_freq/2064,
		half_freq/2065,
		half_freq/2066,
		half_freq/2067,
		half_freq/2068,
		half_freq/2069,
		half_freq/2070,
		half_freq/2071,
		half_freq/2072,
		half_freq/2073,
		half_freq/2074,
		half_freq/2075,
		half_freq/2076,
		half_freq/2077,
		half_freq/2078,
		half_freq/2079,
		half_freq/2080,
		half_freq/2081,
		half_freq/2082,
		half_freq/2083,
		half_freq/2084,
		half_freq/2085,
		half_freq/2086,
		half_freq/2087,
		half_freq/2088,
		half_freq/2089,
		half_freq/2090,
		half_freq/2091,
		half_freq/2092,
		half_freq/2093
	);

	BEGIN
	
	has_space <= '1' when inputs_started = inputs_accepted else '0';
	
	IO_DATA <=
		x"000" & '0' & '0' & '0' & has_space when (SPACE_EN = '1' and IO_WRITE = '0') else
		std_logic_vector(to_unsigned(COMPARE, 16)) when (CS = '1' and IO_WRITE = '0') else
		std_logic_vector(to_unsigned(duration_cycles - duration_cycle_counter, 16)) when (DURATION_EN = '1' and IO_WRITE = '0') else
		(others => 'Z');
	
	PROCESS (CLOCK, RESETN, CS)
	BEGIN
		-- Create a register to store the data sent from SCOMP
		IF (RESETN = '0') THEN
			inputs_accepted <= 0;
			inputs_started <= 0;
			TICKER <= 0;
			
			-- defaults
			next_compare <= 500;
			next_duration_cycles <= -1;
		else
			if rising_edge(CS) and IO_WRITE = '1' then
				if IO_DATA(12 downto 0) <= 2093 then
					next_compare <= conv_integer(IO_DATA(12 downto 0));
				else
					next_compare <= 500;
				end if;
				inputs_accepted <= inputs_accepted + 1;
			end if;
			
			if rising_edge(DURATION_EN) and IO_WRITE = '1' then
				next_duration_cycles <= conv_integer(IO_DATA(15 downto 0));
			end if;
			
			if rising_edge(PAUSE_EN) and IO_WRITE = '1' then
				if IO_DATA = x"0000" then
					PAUSED <= '1';
				else
					PAUSED <= '0';
				end if;
			end if;
			
			if rising_edge(CLOCK) and PAUSED = '0' THEN
				if inputs_accepted > inputs_started then
					-- There is a pending input for us to process
					
					if duration_cycles = -1 then
						-- The currently running frequency has infinite duration; it will not end on its own. Override it immediately.
						COMPARE <= next_compare;
						duration_cycles <= next_duration_cycles;
						duration_cycle_counter <= 0;
						inputs_started <= inputs_started + 1;
						ENABLED <= '1';
						COUNT <= 0;
						TICKER <= 0;
					elsif duration_cycle_counter = duration_cycles then
						-- The currently running frequency has a finite duration and we have completed said duration; switch to the new frequency.
						COMPARE <= next_compare;
						duration_cycles <= next_duration_cycles;
						duration_cycle_counter <= 0;
						inputs_started <= inputs_started + 1;
						ENABLED <= '1';
						COUNT <= 0;
						TICKER <= 0;
					end if;
				elsif duration_cycle_counter = duration_cycles then
					-- We do not have any pending inputs and have reached the end of the current note, so disable it.
					ENABLED <= '0';
				end if;
			
				if ENABLED = '1' then
					if TICKER = 0 and duration_cycles > 0 then
						duration_cycle_counter <= duration_cycle_counter + 1;
					end if;
					TICKER <= TICKER + 1;
				
					IF COUNT < mapping(COMPARE) THEN
						COUNT <= COUNT + 1;
					ELSE
						COUNT <= 0;
						D <= not D and ENABLED;
					END IF;
				else
					D <= '0';
				end if;
			END IF;
		end if;
	END PROCESS;

	SQ <= D;
END a;